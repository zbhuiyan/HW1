module hello_test ();
initial begin
    $display("Hello, CompArch!");
end
endmodule